// AlarmClock_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module AlarmClock_tb (
	);

	wire         alarmclock_inst_clk_bfm_clk_clk;           // AlarmClock_inst_clk_bfm:clk -> [AlarmClock_inst:clk_clk, AlarmClock_inst_reset_bfm:clk]
	wire   [7:0] alarmclock_inst_inputs_bfm_conduit_export; // AlarmClock_inst_inputs_bfm:sig_export -> AlarmClock_inst:inputs_export
	wire  [31:0] alarmclock_inst_leds_export;               // AlarmClock_inst:leds_export -> AlarmClock_inst_leds_bfm:sig_export
	wire         alarmclock_inst_reset_bfm_reset_reset;     // AlarmClock_inst_reset_bfm:reset -> AlarmClock_inst:reset_reset_n

	AlarmClock alarmclock_inst (
		.clk_clk       (alarmclock_inst_clk_bfm_clk_clk),           //    clk.clk
		.inputs_export (alarmclock_inst_inputs_bfm_conduit_export), // inputs.export
		.leds_export   (alarmclock_inst_leds_export),               //   leds.export
		.reset_reset_n (alarmclock_inst_reset_bfm_reset_reset)      //  reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) alarmclock_inst_clk_bfm (
		.clk (alarmclock_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm alarmclock_inst_inputs_bfm (
		.sig_export (alarmclock_inst_inputs_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarmclock_inst_leds_bfm (
		.sig_export (alarmclock_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) alarmclock_inst_reset_bfm (
		.reset (alarmclock_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (alarmclock_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
